module MEMORIA_INSTRUCAO(
	input [11:0] PC,
	output wire [31:0] INSTRUCAO
);
	wire [31:0] memoria[511:0];

	assign memoria[0]={5'd23, 27'd0 }
	assign memoria[1]={5'd23, 27'd0 }
	assign memoria[2]={5'd17, 5'd27, 22'd0 }
	assign memoria[3]={5'd16, 5'd1, 5'd27, 17'd0 }
	assign memoria[4]={5'd17, 5'd27, 22'd13 }
	assign memoria[5]={5'd18, 5'd27, 5'd1, 17'd0 }
	assign memoria[6]={5'd17, 5'd27, 22'd0 }
	assign memoria[7]={5'd16, 5'd2, 5'd27, 17'd0 }
	assign memoria[8]={5'd17, 5'd27, 22'd0 }
	assign memoria[9]={5'd1, 5'd27, 5'd27, 5'd2, 12'd0 }
	assign memoria[10]={5'd16, 5'd3, 5'd27, 17'd0 }
	assign memoria[11]={5'd17, 5'd27, 22'd6 }
	assign memoria[12]={5'd18, 5'd27, 5'd3, 17'd0 }
	assign memoria[13]={5'd17, 5'd27, 22'd0 }
	assign memoria[14]={5'd16, 5'd1, 5'd27, 17'd0 }
	assign memoria[15]={5'd17, 5'd2, 22'd0 }
	assign memoria[16]={5'd1, 5'd3, 5'd1, 5'd2, 12'd0 }
	assign memoria[17]={5'd17, 5'd27, 22'd16 }
	assign memoria[18]={5'd18, 5'd27, 5'd3, 17'd0 }
	assign memoria[19]={5'd23, 27'd0 }
	assign memoria[20]={5'd17, 5'd27, 22'd0 }
	assign memoria[21]={5'd16, 5'd1, 5'd27, 17'd0 }
	assign memoria[22]={5'd17, 5'd27, 22'd0 }
	assign memoria[23]={5'd16, 5'd2, 5'd27, 17'd0 }
	assign memoria[24]={5'd9, 5'd3, 5'd1, 5'd2, 12'd0 }
	assign memoria[25]={5'd11, 5'd3, 5'd0, 17'd3 }
	assign memoria[26]={5'd17, 5'd27, 22'd0 }
	assign memoria[27]={5'd16, 5'd1, 5'd27, 17'd0 }
	assign memoria[28]={5'd17, 5'd27, 22'd0 }
	assign memoria[29]={5'd1, 5'd27, 5'd27, 5'd1, 12'd0 }
	assign memoria[30]={5'd16, 5'd2, 5'd27, 17'd0 }
	assign memoria[31]={5'd17, 5'd27, 22'd0 }
	assign memoria[32]={5'd16, 5'd3, 5'd27, 17'd0 }
	assign memoria[33]={5'd9, 5'd4, 5'd2, 5'd3, 12'd0 }
	assign memoria[34]={5'd11, 5'd4, 5'd0, 17'd4 }
	assign memoria[35]={5'd17, 5'd27, 22'd0 }
	assign memoria[36]={5'd16, 5'd5, 5'd27, 17'd0 }
	assign memoria[37]={5'd17, 5'd27, 22'd0 }
	assign memoria[38]={5'd1, 5'd27, 5'd27, 5'd5, 12'd0 }
	assign memoria[39]={5'd16, 5'd6, 5'd27, 17'd0 }
	assign memoria[40]={5'd17, 5'd27, 22'd6 }
	assign memoria[41]={5'd18, 5'd27, 5'd6, 17'd0 }
	assign memoria[42]={5'd17, 5'd27, 22'd0 }
	assign memoria[43]={5'd16, 5'd7, 5'd27, 17'd0 }
	assign memoria[44]={5'd17, 5'd27, 22'd13 }
	assign memoria[45]={5'd18, 5'd27, 5'd7, 17'd0 }
	assign memoria[46]={5'd23, 27'd0 }
	assign memoria[47]={5'd17, 5'd27, 22'd0 }
	assign memoria[48]={5'd16, 5'd8, 5'd27, 17'd0 }
	assign memoria[49]={5'd17, 5'd9, 22'd0 }
	assign memoria[50]={5'd1, 5'd10, 5'd8, 5'd9, 12'd0 }
	assign memoria[51]={5'd17, 5'd27, 22'd16 }
	assign memoria[52]={5'd18, 5'd27, 5'd10, 17'd0 }
	assign memoria[53]={5'd13, 27'd19 }
	assign memoria[54]={5'd23, 27'd0 }
	assign memoria[55]={5'd17, 5'd27, 22'd0 }
	assign memoria[56]={5'd16, 5'd11, 5'd27, 17'd0 }
	assign memoria[57]={5'd19, 5'd28, 5'd11, 17'd0 }
	assign memoria[58]={5'd14, 5'd31, 22'd0 }
	assign memoria[59]={5'd14, 5'd31, 22'd0 }
	assign memoria[60]={5'd23, 27'd0 }
	assign memoria[61]={5'd17, 5'd27, 22'd0 }
	assign memoria[62]={5'd16, 5'd12, 5'd27, 17'd0 }
	assign memoria[63]={5'd17, 5'd27, 22'd16 }
	assign memoria[64]={5'd18, 5'd27, 5'd12, 17'd0 }
	assign memoria[65]={5'd23, 27'd0 }
	assign memoria[66]={5'd17, 5'd27, 22'd0 }
	assign memoria[67]={5'd16, 5'd13, 5'd27, 17'd0 }
	assign memoria[68]={5'd17, 5'd14, 22'd0 }
	assign memoria[69]={5'd2, 5'd15, 5'd13, 5'd14, 12'd0 }
	assign memoria[70]={5'd17, 5'd27, 22'd0 }
	assign memoria[71]={5'd16, 5'd16, 5'd27, 17'd0 }
	assign memoria[72]={5'd9, 5'd17, 5'd16, 5'd15, 12'd0 }
	assign memoria[73]={5'd11, 5'd17, 5'd0, 17'd7 }
	assign memoria[74]={5'd17, 5'd27, 22'd0 }
	assign memoria[75]={5'd16, 5'd18, 5'd27, 17'd0 }
	assign memoria[76]={5'd19, 5'd22, 5'd18, 17'd0 }
	assign memoria[77]={5'd17, 5'd27, 22'd0 }
	assign memoria[78]={5'd16, 5'd19, 5'd27, 17'd0 }
	assign memoria[79]={5'd19, 5'd23, 5'd19, 17'd0 }
	assign memoria[80]={5'd17, 5'd27, 22'd0 }
	assign memoria[81]={5'd16, 5'd20, 5'd27, 17'd0 }
	assign memoria[82]={5'd19, 5'd24, 5'd20, 17'd0 }
	assign memoria[83]={5'd15, 27'd0 }
	assign memoria[84]={5'd19, 5'd21, 5'd28, 17'd0 }
	assign memoria[85]={5'd17, 5'd27, 22'd13 }
	assign memoria[86]={5'd18, 5'd27, 5'd21, 17'd0 }
	assign memoria[87]={5'd17, 5'd27, 22'd0 }
	assign memoria[88]={5'd16, 5'd22, 5'd27, 17'd0 }
	assign memoria[89]={5'd17, 5'd27, 22'd0 }
	assign memoria[90]={5'd1, 5'd27, 5'd27, 5'd22, 12'd0 }
	assign memoria[91]={5'd16, 5'd23, 5'd27, 17'd0 }
	assign memoria[92]={5'd17, 5'd27, 22'd14 }
	assign memoria[93]={5'd18, 5'd27, 5'd23, 17'd0 }
	assign memoria[94]={5'd17, 5'd27, 22'd0 }
	assign memoria[95]={5'd16, 5'd24, 5'd27, 17'd0 }
	assign memoria[96]={5'd17, 5'd27, 22'd0 }
	assign memoria[97]={5'd1, 5'd27, 5'd27, 5'd24, 12'd0 }
	assign memoria[98]={5'd16, 5'd25, 5'd27, 17'd0 }
	assign memoria[99]={5'd17, 5'd27, 22'd0 }
	assign memoria[100]={5'd16, 5'd26, 5'd27, 17'd0 }
	assign memoria[101]={5'd17, 5'd27, 22'd9 }
	assign memoria[102]={5'd1, 5'd27, 5'd27, 5'd26, 12'd0 }
	assign memoria[103]={5'd18, 5'd27, 5'd25, 17'd0 }
	assign memoria[104]={5'd17, 5'd27, 22'd0 }
	assign memoria[105]={5'd16, 5'd27, 5'd27, 17'd0 }
	assign memoria[106]={5'd17, 5'd27, 22'd0 }
	assign memoria[107]={5'd16, 5'd28, 5'd27, 17'd0 }
	assign memoria[108]={5'd17, 5'd27, 22'd9 }
	assign memoria[109]={5'd1, 5'd27, 5'd27, 5'd28, 12'd0 }
	assign memoria[110]={5'd18, 5'd27, 5'd27, 17'd0 }
	assign memoria[111]={5'd17, 5'd27, 22'd0 }
	assign memoria[112]={5'd16, 5'd29, 5'd27, 17'd0 }
	assign memoria[113]={5'd17, 5'd30, 22'd0 }
	assign memoria[114]={5'd1, 5'd31, 5'd29, 5'd30, 12'd0 }
	assign memoria[115]={5'd17, 5'd27, 22'd16 }
	assign memoria[116]={5'd18, 5'd27, 5'd31, 17'd0 }
	assign memoria[117]={5'd13, 27'd65 }
	assign memoria[118]={5'd23, 27'd0 }
	assign memoria[119]={5'd14, 5'd31, 22'd0 }
	assign memoria[120]={5'd23, 27'd0 }
	assign memoria[121]={5'd17, 5'd32, 22'd0 }
	assign memoria[122]={5'd17, 5'd27, 22'd16 }
	assign memoria[123]={5'd18, 5'd27, 5'd32, 17'd0 }
	assign memoria[124]={5'd23, 27'd0 }
	assign memoria[125]={5'd17, 5'd27, 22'd0 }
	assign memoria[126]={5'd16, 5'd33, 5'd27, 17'd0 }
	assign memoria[127]={5'd17, 5'd34, 22'd0 }
	assign memoria[128]={5'd9, 5'd35, 5'd33, 5'd34, 12'd0 }
	assign memoria[129]={5'd11, 5'd35, 5'd0, 17'd10 }
	assign memoria[130]={5'd20, 27'd0 }
	assign memoria[131]={5'd19, 5'd36, 5'd30, 17'd0 }
	assign memoria[132]={5'd17, 5'd27, 22'd0 }
	assign memoria[133]={5'd16, 5'd37, 5'd27, 17'd0 }
	assign memoria[134]={5'd17, 5'd27, 22'd0 }
	assign memoria[135]={5'd1, 5'd27, 5'd27, 5'd37, 12'd0 }
	assign memoria[136]={5'd18, 5'd27, 5'd36, 17'd0 }
	assign memoria[137]={5'd17, 5'd27, 22'd0 }
	assign memoria[138]={5'd16, 5'd38, 5'd27, 17'd0 }
	assign memoria[139]={5'd17, 5'd39, 22'd0 }
	assign memoria[140]={5'd1, 5'd40, 5'd38, 5'd39, 12'd0 }
	assign memoria[141]={5'd17, 5'd27, 22'd16 }
	assign memoria[142]={5'd18, 5'd27, 5'd40, 17'd0 }
	assign memoria[143]={5'd13, 27'd124 }
	assign memoria[144]={5'd23, 27'd0 }
	assign memoria[145]={5'd17, 5'd27, 22'd0 }
	assign memoria[146]={5'd16, 5'd41, 5'd27, 17'd0 }
	assign memoria[147]={5'd19, 5'd25, 5'd41, 17'd0 }
	assign memoria[148]={5'd17, 5'd42, 22'd0 }
	assign memoria[149]={5'd19, 5'd26, 5'd42, 17'd0 }
	assign memoria[150]={5'd17, 5'd43, 22'd0 }
	assign memoria[151]={5'd19, 5'd27, 5'd43, 17'd0 }
	assign memoria[152]={5'd15, 27'd0 }
	assign memoria[153]={5'd17, 5'd44, 22'd0 }
	assign memoria[154]={5'd17, 5'd27, 22'd16 }
	assign memoria[155]={5'd18, 5'd27, 5'd44, 17'd0 }
	assign memoria[156]={5'd23, 27'd0 }
	assign memoria[157]={5'd17, 5'd27, 22'd0 }
	assign memoria[158]={5'd16, 5'd45, 5'd27, 17'd0 }
	assign memoria[159]={5'd17, 5'd46, 22'd0 }
	assign memoria[160]={5'd9, 5'd47, 5'd45, 5'd46, 12'd0 }
	assign memoria[161]={5'd11, 5'd47, 5'd0, 17'd12 }
	assign memoria[162]={5'd17, 5'd27, 22'd0 }
	assign memoria[163]={5'd16, 5'd48, 5'd27, 17'd0 }
	assign memoria[164]={5'd17, 5'd27, 22'd0 }
	assign memoria[165]={5'd1, 5'd27, 5'd27, 5'd48, 12'd0 }
	assign memoria[166]={5'd16, 5'd49, 5'd27, 17'd0 }
	assign memoria[167]={5'd19, 5'd28, 5'd49, 17'd0 }
	assign memoria[168]={5'd24, 5'd22, 22'd0 }
	assign memoria[169]={5'd17, 5'd27, 22'd0 }
	assign memoria[170]={5'd16, 5'd50, 5'd27, 17'd0 }
	assign memoria[171]={5'd17, 5'd51, 22'd0 }
	assign memoria[172]={5'd1, 5'd52, 5'd50, 5'd51, 12'd0 }
	assign memoria[173]={5'd17, 5'd27, 22'd16 }
	assign memoria[174]={5'd18, 5'd27, 5'd52, 17'd0 }
	assign memoria[175]={5'd13, 27'd156 }
	assign memoria[176]={5'd23, 27'd0 }
	assign memoria[177]={5'd21, 27'd0 }

	assign INSTRUCAO = memoria [PC]; 

endmodule
